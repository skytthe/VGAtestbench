library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity vga_generator is
	port (
		clk_i : in std_logic
	);
end entity vga_generator;

architecture Behavioral of vga_generator is
	
begin
	
end architecture Behavioral;

