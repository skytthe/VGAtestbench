library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity vga_sampler is
	port (
		clk_i : in std_logic
	);
end entity vga_sampler;

architecture Behavioral of vga_sampler is

	signal tk : std_logic;
	
	
begin


	
end architecture Behavioral;
